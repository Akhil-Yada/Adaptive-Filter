  module d2(y,x,w1,w,t,r,clk);
  output [9:0]y;
  input [7:0]x;
  input [9:0]w;
  input w1,t,r,clk;
  wire c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,s1,s2,s3,s4,s5,s6,s7,s8,s9,s10;
  wire a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,b1,b2,b3,b4,b5,b6,b7,b8,b9,b10;
  assign y={s1,s2,s3,s4,s5,s6,s7,s8,s9,s10};
  ///////////////////////////////////////////////////////////////////////////////////////
  assign a1=(s1&t);
  assign a2=(x[7]&~t)|(s2&t);
  assign a3=(x[6]&~t)|(s3&t);
  assign a4=(x[5]&~t)|(s4&t);
  assign a5=(x[4]&~t)|(s5&t);
  assign a6=(x[3]&~t)|(s6&t);
  assign a7=(x[2]&~t)|(s7&t);
  assign a8=(x[1]&~t)|(s8&t);
  assign a9=(x[0]&~t)|(s9&t);
  //////////////////////////////////////////////////////////////////////////////////////
  assign b1=(c1&t)|(w1&~t);
  assign b2=(c2&t)|(w1&~t);
  assign b3=(c3&t)|(w1&~t);
  assign b4=(c4&t)|(w1&~t);
  assign b5=(c5&t)|(w1&~t);
  assign b6=(c6&t)|(w1&~t);
  assign b7=(c7&t)|(w1&~t);
  assign b8=(c8&t)|(w1&~t);
  assign b9=(c9&t)|(w1&~t);
  assign b10=(c10&t)|(w1&~t);
  //////////////////////////////////////////////////////////////////////////////////////
  csa cs1(s1,c1,w[9],a1,b1,r,clk);
  csa cs2(s2,c2,w[8],a1,b2,r,clk);
  csa cs3(s3,c3,w[7],a2,b3,r,clk);
  csa cs4(s4,c4,w[6],a3,b4,r,clk);
  csa cs5(s5,c5,w[5],a4,b5,r,clk);
  csa cs6(s6,c6,w[4],a5,b6,r,clk);
  csa cs7(s7,c7,w[3],a6,b7,r,clk);
  csa cs8(s8,c8,w[2],a7,b8,r,clk);
  csa cs9(s9,c9,w[3],a8,b9,r,clk);
  csa cs10(s10,c10,w[2],a9,b10,r,clk);
endmodule

module test_design2();
reg [3:0]a;
reg r,clk;
d2 testd2(a,r,clk);
initial
begin
r=0;
#10;
r=1;
#10;
clk=0;
#80;
//////////////////////////////////////////////////
a=4'b0111;
#50;
clk=1;
#50;
////////////////////////////////////////////
clk=0;
#10;
a=4'b1010;
#50
clk=1;
#40;
////////////////////////////////////////////
clk=0;
#10;
a=4'b1101;
#50
clk=1;
#40;
////////////////////////////////////////////
clk=0;
#10;
a=4'b1011;
#50
clk=1;
#40;
////////////////////////////////////////////
clk=0;
#10;
a=4'b0000;
#50
clk=1;
#40;
////////////////////////////////////////////
clk=0;
#10;
a=4'b0000;
#50
clk=1;
#40;
////////////////////////////////////////////
clk=0;
#10;
a=4'b0000;
#50
clk=1;
#40;
////////////////////////////////////////////
end
endmodule