module iptb(A2,A3,A4,A5,A6,A7,A8,A9,A10,A11,A12,A13,A14,A15,A16,x1,x2,x3,r,clk);
input [7:0]x1,x2,x3;
input r,clk;
output [9:0]A2,A3,A4,A5,A6,A7,A8,A9,A10,A11,A12,A13,A14,A15,A16;
wire [7:0]x4;
wire [8:0]a,b,c,d,e,f;
assign a={x1[7],x1}+{x2[7],x2};//x(n)+x(n-1)
assign b={x1[7],x1}+{x3[7],x3};//x(n)+x(n-2)
assign c={x1[7],x1}+{x4[7],x4};//x(n)+x(n-3)
assign A15={x1[7],x1[7],x1}+{d[8],d};//x(n)+x(n-1)+x(n-2)
assign A12={x1[7],x1[7],x1}+{f[8],f};//x(n)+x(n-2)+x(n-3)
assign A14={x1[7],x1[7],x1}+{e[8],e};//x(n)+x(n-1)+x(n-3)
assign A16={x1[7],x1[7],x1}+A8;//x(n)+x(n-1)+x(n-2)+x(n-3)
assign A13={a[8],a};
assign A11={b[8],b};
assign A10={c[8],c};
assign A7={d[8],d};
assign A6={e[8],e};
assign A4={f[8],f};
assign A9={x1[7],x1[7],x1};//x(n)
assign A5={x2[7],x2[7],x2};//x(n-1)
assign A3={x3[7],x3[7],x3};//x(n-2)
assign A2={x4[7],x4[7],x4};//x(n-3)
Dffp df1[7:0](x4,x3,r,clk); 
Dffp df2[8:0](d,a,r,clk);//x(n-1)+x(n-2)
Dffp df3[8:0](f,d,r,clk);//x(n-2)+x(n-3)
Dffp df4[8:0](e,b,r,clk);//x(n-1)+x(n-3)
Dffp df5[9:0](A8,A15,r,clk);//x(n-1)+x(n-2)+x(n-3)
endmodule