 module cc(cc1,cc2,w1,x1,a,b,s0,s1,s2);
 input [7:0]w1,x1;
 input a,b,s0,s1,s2;
 output cc1,cc2;
 wire c0,c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16;
 wire [7:0]w,x;
 xor xr1[7:0](w,w1,b);
 xor xr2[7:0](x,x1,a);
 assign c0=(w[0]&(x[0]|a|b)|x[0]&(a|b)|a&b)&~c1;
 assign c1=w[0]&x[0]&a&b;
 assign c2=s0&c1;
 assign c3=c1&~s0;
 //////////////////////////////////////////////////////////////////////////////////////
 assign c4=s0&(w[1]&(x[1]|c0)|x[1]&c0)|~s0&c0; 
 //////////////////////////////////////////////////////////////////////////////////////
 assign c5=s1&((w[2]&(x[2]|c4|c2)|x[2]&(c4|c2)|c4&c2)&~c6);
 assign c6=s1&((w[2]&x[2]&c4&c2))|~s1&c4;
 assign c7=s1&((w[3]&(x[3]|c5|c3)|x[3]&(c5|c3)|c5&c3)&~c8)|~s1&c2;
 assign c8=s1&(w[3]&x[3]&c3&c5)|~s1&c3;
 /////////////////////////////////////////////////////////////////////////////////////
 assign c9=(w[4]&(x[4]|c6|c7)|x[4]&(c6|c7)|c6&c7)&~c10;
 assign c10=w[4]&x[4]&c6&c7;
 assign c11=(w[5]&(x[5]|c9|c8)|x[5]&(c9|c8)|c9&c8)&~c12;
 assign c12=w[5]&x[5]&c9&c8;
 assign c13=(w[6]&(x[6]|c11|c10)|x[6]&(c11|c10)|c11&c10)&~c14;
 assign c14=w[6]&x[6]&c11&c10;
 assign c15=(w[7]&(x[7]|c12|c13)|x[7]&(c12|c13)|c12&c13)&~c16;
 assign c16=w[7]&x[7]&c12&c13;
 ///////////////////////////////////////////////////////////////////////////////////////
 assign cc1=~s2&(c6|c8)|s2&(c14|c16);
 assign cc2=~s2&(c7|c8)|s2&(c15|c16);
endmodule
