module bsmb(o,w,s0,s1,s2,x);
 input s0,s1,s2,x;
 input [9:0]w;
 output [9:0]o;
 wire [9:0]l1,l2,l3;
 and r1_1(l1[9],w[9],x);
 and r1_2(l1[8],w[8],x);
 and r1_3(l1[7],w[7],x);
 and r1_4(l1[6],w[6],x);
 and r1_5(l1[5],w[5],x);
 and r1_6(l1[4],w[4],x);
 and r1_7(l1[3],w[3],x);
 and r1_8(l1[2],w[2],x);
 and r1_9(l1[1],w[1],x);
 and r1_10(l1[0],w[0],x);
 ///////////////////////////////////////////////////////////////
 Mux2_1 r2_1(l2[9],l1[9],l1[9],s0);
 Mux2_1 r2_2(l2[8],l1[8],l1[9],s0);
 Mux2_1 r2_3(l2[7],l1[7],l1[8],s0);
 Mux2_1 r2_4(l2[6],l1[6],l1[7],s0);
 Mux2_1 r2_5(l2[5],l1[5],l1[6],s0);
 Mux2_1 r2_6(l2[4],l1[4],l1[5],s0);
 Mux2_1 r2_7(l2[3],l1[3],l1[4],s0); 
 Mux2_1 r2_8(l2[2],l1[2],l1[3],s0);
 Mux2_1 r2_9(l2[1],l1[1],l1[2],s0); 
 Mux2_1 r2_10(l2[0],l1[0],l1[1],s0);
 ///////////////////////////////////////////////////////////////
 Mux2_1 r3_1(l3[9],l2[9],l2[9],s1);
 Mux2_1 r3_2(l3[8],l2[8],l2[9],s1);
 Mux2_1 r3_3(l3[7],l2[7],l2[9],s1);
 Mux2_1 r3_4(l3[6],l2[6],l2[8],s1);
 Mux2_1 r3_5(l3[5],l2[5],l2[7],s1);
 Mux2_1 r3_6(l3[4],l2[4],l2[6],s1);
 Mux2_1 r3_7(l3[3],l2[3],l2[5],s1); 
 Mux2_1 r3_8(l3[2],l2[2],l2[4],s1);
 Mux2_1 r3_9(l3[1],l2[1],l2[3],s1); 
 Mux2_1 r3_10(l3[0],l2[0],l2[2],s1);
 /////////////////////////////////////////////////////////////////
 Mux2_1 r4_1(o[9],l3[9],l3[9],s2);
 Mux2_1 r4_2(o[8],l3[8],l3[9],s2);
 Mux2_1 r4_3(o[7],l3[7],l2[9],s2);
 Mux2_1 r4_4(o[6],l3[6],l3[9],s2);
 Mux2_1 r4_5(o[5],l3[5],l3[9],s2);
 Mux2_1 r4_6(o[4],l3[4],l3[8],s2);
 Mux2_1 r4_7(o[3],l3[3],l3[7],s2); 
 Mux2_1 r4_8(o[2],l3[2],l3[6],s2);
 Mux2_1 r4_9(o[1],l3[1],l3[5],s2); 
 Mux2_1 r4_10(o[0],l3[0],l3[4],s2);
 endmodule
