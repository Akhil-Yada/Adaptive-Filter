 module iptm(x10,A1,A2,A3,A4,x,x_,r,clk);
 input [7:0]x,x_;
 input r,clk;
 output [9:0]A1,A2,A3,A4,x10;
 wire [7:0]x_,xn_,x;
 wire [8:0]R1o,R1i,R2o,R2i;
 wire [9:0]R3i,R4i,R5i,R6i;
 wire [8:0]c1,c2;
 wire [9:0]r1o,r2o;
 
 Dffp R1[8:0](R1o,R1i,r,clk);
 Dffp R2[8:0](R2o,R2i,r,clk);
 Dffp R3[9:0](A1,R3i,r,clk);
 Dffp R4[9:0](A2,R4i,r,clk);
 Dffp R5[9:0](A3,R5i,r,clk);
 Dffp R6[9:0](A4,R6i,r,clk);
 /////////////////////////////////////////////////////////////////////////////////////////////////////
 FA f1(R1i[0],c1[0],x[0],x_[0],1'b0);
 FA f2(R1i[1],c1[1],x[1],x_[1],c1[0]);
 FA f3(R1i[2],c1[2],x[2],x_[2],c1[1]);
 FA f4(R1i[3],c1[3],x[3],x_[3],c1[2]);
 FA f5(R1i[4],c1[4],x[4],x_[4],c1[3]);
 FA f6(R1i[5],c1[5],x[5],x_[5],c1[4]);
 FA f7(R1i[6],c1[6],x[6],x_[6],c1[5]);
 FA f8(R1i[7],c1[7],x[7],x_[7],c1[6]);
 FA f9(R1i[8],c1[8],x[7],x_[7],c1[7]);
 ////////////////////////////////////////////////////////////////////////////////////////////////////
 not n[7:0](xn_,x_);
 FA q1(R2i[0],c2[0],x[0],xn_[0],1'b1);
 FA q2(R2i[1],c2[1],x[1],xn_[1],c2[0]);
 FA q3(R2i[2],c2[2],x[2],xn_[2],c2[1]);
 FA q4(R2i[3],c2[3],x[3],xn_[3],c2[2]);
 FA q5(R2i[4],c2[4],x[4],xn_[4],c2[3]);
 FA q6(R2i[5],c2[5],x[5],xn_[5],c2[4]);
 FA q7(R2i[6],c2[6],x[6],xn_[6],c2[5]);
 FA q8(R2i[7],c2[7],x[7],xn_[7],c2[6]);
 FA q9(R2i[8],c2[8],x[7],xn_[7],c2[7]);
 /////////////////////////////////////////////////////////////////////////////////////////////////////
 assign x10={x[7],x[7],x};
 assign r1o={R1o[8],R1o};
 assign r2o={R2o[8],R2o};
 add10 a1(R3i,x10,r1o);
 sub10 s1(R4i,x10,r1o);
 add10 a2(R5i,x10,r2o);
 sub10 s2(R6i,x10,r2o);
 endmodule