module DA11(sum,carry,t,x1,x2,x3,x4,w1,w2,w3,w4,w5,w6,w7,w8,r,clk);
output [10:0]sum,carry;
input [5:0]t;
input [7:0]x1,x2,x3,x4;
input [9:0]w1,w2,w3,w4,w5,w6,w7,w8;
input r,clk;
wire t5,t6,t_,z;
wire a,a_,b,b_,c,c_,d,d_,e,e_,f,f_,g,g_,h,h_;
wire [9:0]l1,l2,l1_,l2_,lx1,lx2,w;
wire [7:0]x1_;
assign {t6,t5,z4,z3,z2,z1}=t;
assign t_=~t6;
assign z=~(t5|t6);
///////////////////////////////////////////////////////////////////////////////////////////////////
assign a=(z1&x1[0])|(z2&x1[2])|(z3&x1[4])|(z4&x1[6]);
assign b=(z2&x2[0])|(z2&x2[2])|(z3&x2[4])|(z4&x2[6]);
assign c=(z3&x3[0])|(z2&x3[2])|(z3&x3[4])|(z4&x3[6]);
assign d=(z4&x4[0])|(z2&x4[2])|(z3&x4[4])|(z4&x4[6]);  
///////////////////////////////////////////////////////////////////////////////////////////////////
assign e=(z1&x1[1])|(z2&x1[3])|(z3&x1[5])|(z4&~x1[7]);
assign f=(z2&x2[1])|(z2&x2[3])|(z3&x2[5])|(z4&~x2[7]);
assign g=(z3&x3[1])|(z2&x3[3])|(z3&x3[5])|(z4&~x3[7]);
assign h=(z4&x4[1])|(z2&x4[3])|(z3&x4[5])|(z4&~x4[7]); 
//////////////////////////////////////////////////////////////////////////////////////////////////
assign x1_={x1[7],~x1[6],~x1[5],~x1[4],~x1[3],~x1[2],~x1[1],~x1[0]};
not nw[9:0](w,w1);
not (a_,a);
not (e_,e);
xor (b_,b,a);
xor (c_,c,a);
xor (d_,d,a);
xor (f_,f,e);
xor (g_,g,e);
xor (h_,h,e);
mux8_18 m1(l1,w1,w2,w3,w4,w5,w6,w7,w8,b_,c_,d_);
mux8_18 m2(l2,w1,w2,w3,w4,w5,w6,w7,w8,f_,g_,h_);
xor xr1[9:0](lx1,l1,a_);
xor xr2[9:0](lx2,l2,e_);
and a1[9:0](l1_,lx1,z);
and a2[9:0](l2_,lx2,z);
/////////////////////////////////////////////////////////////////////////////////////////////////
d1 mac(sum,carry,x1_,w,l2_,l1_,t_,r,clk);
endmodule
